module Instruction_Memory(
    input clk, rst,
    input[31:0] address, 
    output reg[31:0] instruction
);
    reg[7:0] data [0:1023];
    always @(*) begin
        if (rst)
        begin
            instruction <= 32'b0;
            {data[0], data[1], data[2], data[3]} =      32'b1110_00_1_1101_0_0000_0000_000000010100; //MOV R0 ,#20 //R0 = 20
            {data[4], data[5], data[6], data[7]} =      32'b1110_00_1_1101_0_0000_0001_101000000001; //MOV R1 ,#4096 //R1 = 4096
            {data[8], data[9], data[10], data[11]} =    32'b1110_00_1_1101_0_0000_0010_000100000011; //MOV R2 ,#0xC0000000 //R2 = -1073741824
            {data[12], data[13], data[14], data[15]} =  32'b1110_00_0_0100_1_0010_0011_000000000010; //ADDS R3 ,R2,R2 //R3 = -2147483648
            {data[16], data[17], data[18], data[19]} =  32'b1110_00_0_0101_0_0000_0100_000000000000; //ADC R4 ,R0,R0 //R4 = 41
            {data[20], data[21], data[22], data[23]} =  32'b1110_00_0_0010_0_0100_0101_000100000100; //SUB R5 ,R4,R4,LSL #2 //R5 = -123
            {data[24], data[25], data[26], data[27]} =  32'b1110_00_0_0110_0_0000_0110_000010100000; //SBC R6 ,R0,R0,LSR #1 //R6 = -10
            {data[28], data[29], data[30], data[31]} =  32'b1110_00_0_1100_0_0101_0111_000101000010; //ORR R7 ,R5,R2,ASR #2 //R7 = -123
            {data[32], data[33], data[34], data[35]} =  32'b1110_00_0_0000_0_0111_1000_000000000011; //AND R8 ,R7,R3 //R8 = -2147483648
            {data[36], data[37], data[38], data[39]} =  32'b1110_00_0_1111_0_0000_1001_000000000110; //MVN R9 ,R6 //R9 = 10
            {data[40], data[41], data[42], data[43]} =  32'b1110_00_0_0001_0_0100_1010_000000000101; //EOR R10,R4,R5 //R10 = -84
            {data[44], data[45], data[46], data[47]} =  32'b1110_00_0_1010_1_1000_0000_000000000110; //CMP R8 ,R6
            {data[48], data[49], data[50], data[51]} =  32'b0001_00_0_0100_0_0001_0001_000000000001; //ADDNE R1 ,R1,R1 //R1 = 8192
            {data[52], data[53], data[54], data[55]} =  32'b1110_00_0_1000_1_1001_0000_000000001000; //TST R9 ,R8
            {data[56], data[57], data[58], data[59]} =  32'b0000_00_0_0100_0_0010_0010_000000000010; //ADDEQ R2 ,R2,R2 //R2 = -1073741824
            {data[60], data[61], data[62], data[63]} =  32'b1110_00_1_1101_0_0000_0000_101100000001; //MOV R0 ,#1024 //R0 = 1024
            {data[64], data[65], data[66], data[67]} =  32'b1110_01_0_0100_0_0000_0001_000000000000; //STR R1 ,[R0],#0 //MEM[1024] = 8192
            {data[68], data[69], data[70], data[71]} =  32'b1110_01_0_0100_1_0000_1011_000000000000; //LDR R11,[R0],#0 //R11 = 8192
        end
        else
        begin
            instruction <= {data[address],data[address+1],data[address+2],data[address+3]};
        end
    end
    
endmodule